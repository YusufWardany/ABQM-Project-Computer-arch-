module Rom(
input clk, 
input reset, 
input [4:0] address,
           
output reg [7:0] data_out);
           
    always @(posedge clk or posedge reset) begin
if(reset)
begin
data_out = 8'b00000000;
end
else
begin
        case(address)
            5'b01000 : data_out = 8'b00000000;
            5'b01001 : data_out = 8'b00000011;
            5'b01010 : data_out = 8'b00000110;
            5'b01011 : data_out = 8'b00001001;
            5'b01100 : data_out = 8'b00010010;
            5'b01101 : data_out = 8'b00010101;
            5'b01110 : data_out = 8'b00011000;
            5'b01111 : data_out = 8'b00100001;
            5'b10000 : data_out = 8'b00000000;
            5'b10001 : data_out = 8'b00000011;
            5'b10010 : data_out = 8'b00000100;
            5'b10011 : data_out = 8'b00000110;
            5'b10100 : data_out = 8'b00000111;
            5'b10101 : data_out = 8'b00001001;
            5'b10110 : data_out = 8'b00010000;
            5'b10111 : data_out = 8'b00010010;
            5'b11000 : data_out = 8'b00000000;
            5'b11001 : data_out = 8'b00000011;
            5'b11010 : data_out = 8'b00000100;
            5'b11011 : data_out = 8'b00000101;
            5'b11100 : data_out = 8'b00000110;
            5'b11101 : data_out = 8'b00000111;
            5'b11110 : data_out = 8'b00001000;
            5'b11111: data_out = 8'b00001001;
            default: data_out = 8'b00000000;
        endcase
end
    end
    
endmodule

